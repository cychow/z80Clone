module z80_alu(

);

endmodule
