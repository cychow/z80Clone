

module z80_regs(
    input clk,
    input rst_n,
    inout [7:0] data
    
);

// reg [7:0] 
/*
always @(posedge clk, negedge rst_n) begin
    

end
*/
endmodule
