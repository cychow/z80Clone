module z80_decode (

);


endmodule
