// z80_decode: instruction decoding

module z80_decode (

);


endmodule
