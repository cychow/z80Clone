module z80_alu(
    input clk,
    input rst_n,
    inout [7:0] data
);



endmodule
