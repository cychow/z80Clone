

module z80_regs(
    input clk,
    input rst_n,
    input [7:0] data,
    
);

always @(posedge clk, negedge rst_n) begin
    

end

endmodule
